// TODO

`default_nettype none

module TODO #(
        parameter TODO = TODO
    ) (
        input wire clk,
        input wire rst,

        input wire TODO,
        output logic TODO
    );

endmodule

`default_nettype wire
